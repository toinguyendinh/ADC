magic
tech sky130A
timestamp 1692049728
<< error_s >>
rect 600 1150 627 1550
rect 2050 1150 2077 1550
rect 1050 800 1077 1150
rect 2500 800 2527 1150
<< nwell >>
rect 1300 800 1450 820
rect 2750 800 2900 820
<< pwell >>
rect 1300 630 1450 650
rect 2750 630 2900 650
<< poly >>
rect 100 630 250 820
rect 550 750 600 770
rect 450 700 600 750
rect 550 280 600 700
rect 950 750 1000 1170
rect 950 700 1100 750
rect 950 680 1000 700
rect 1300 630 1450 820
rect 1550 630 1700 820
rect 2000 750 2050 770
rect 1900 700 2050 750
rect 2000 280 2050 700
rect 2400 750 2450 1170
rect 2400 700 2550 750
rect 2400 680 2450 700
rect 2750 630 2900 820
<< locali >>
rect 70 1442 100 1550
rect 300 1150 450 1200
rect 520 1112 550 1550
rect 1450 1442 1480 1550
rect 1520 1442 1550 1550
rect 1800 1350 1900 1400
rect 120 670 230 780
rect 450 750 480 838
rect 620 750 650 1188
rect 1970 1112 2000 1550
rect 2900 1442 2930 1550
rect 450 700 650 750
rect 450 612 480 700
rect 620 662 650 700
rect 900 750 930 788
rect 1070 750 1100 838
rect 900 700 1100 750
rect 900 262 930 700
rect 1070 612 1100 700
rect 1320 670 1430 780
rect 1570 670 1680 780
rect 1900 750 1930 838
rect 2070 750 2100 1188
rect 1900 700 2100 750
rect 1900 612 1930 700
rect 2070 662 2100 700
rect 2350 750 2380 788
rect 2520 750 2550 838
rect 2350 700 2550 750
rect 70 -100 100 8
rect 1000 -100 1030 338
rect 2350 262 2380 700
rect 2520 612 2550 700
rect 2770 670 2880 780
rect 1450 -100 1480 8
rect 1520 -100 1550 8
rect 2450 -100 2480 338
rect 2550 50 2650 100
rect 2900 -100 2930 8
<< metal1 >>
rect 300 1050 350 1200
rect 50 1000 200 1050
rect 300 1000 1650 1050
rect 150 780 200 1000
rect 1600 780 1650 1000
rect 120 670 230 780
rect 1320 670 1430 780
rect 1570 670 1680 780
rect 2770 670 2880 780
rect 1350 450 1400 670
rect 2800 500 2850 670
rect 1700 450 2850 500
rect 1700 350 1750 450
rect 1250 300 1750 350
use nfet_12  nfet_12_0
timestamp 1692025688
transform 1 0 2450 0 1 110
box 50 -140 500 540
use nfet_12  nfet_12_1
timestamp 1692025688
transform 1 0 1450 0 1 110
box 50 -140 500 540
use nfet_12  nfet_12_2
timestamp 1692025688
transform 1 0 0 0 1 110
box 50 -140 500 540
use nfet_12  nfet_12_3
timestamp 1692025688
transform 1 0 1000 0 1 110
box 50 -140 500 540
use nfet_34  nfet_34_0
timestamp 1692022408
transform 1 0 2100 0 1 340
box -50 -40 400 360
use nfet_34  nfet_34_1
timestamp 1692022408
transform 1 0 2000 0 1 -60
box -50 -40 400 360
use nfet_34  nfet_34_2
timestamp 1692022408
transform 1 0 550 0 1 -60
box -50 -40 400 360
use nfet_34  nfet_34_3
timestamp 1692022408
transform 1 0 650 0 1 340
box -50 -40 400 360
use pfet_12  pfet_12_0
timestamp 1692027968
transform 1 0 2500 0 1 800
box 0 0 450 680
use pfet_12  pfet_12_1
timestamp 1692027968
transform 1 0 1500 0 1 800
box 0 0 450 680
use pfet_12  pfet_12_2
timestamp 1692027968
transform 1 0 50 0 1 800
box 0 0 450 680
use pfet_12  pfet_12_3
timestamp 1692027968
transform 1 0 1050 0 1 800
box 0 0 450 680
use pfet_34  pfet_34_0
timestamp 1692022863
transform 1 0 2100 0 1 1190
box -50 -40 400 360
use pfet_34  pfet_34_1
timestamp 1692022863
transform 1 0 2000 0 1 790
box -50 -40 400 360
use pfet_34  pfet_34_2
timestamp 1692022863
transform 1 0 550 0 1 790
box -50 -40 400 360
use pfet_34  pfet_34_3
timestamp 1692022863
transform 1 0 650 0 1 1190
box -50 -40 400 360
<< end >>
