magic
tech sky130A
timestamp 1692025688
<< pwell >>
rect 50 -140 500 540
<< nmos >>
rect 100 -100 450 500
<< ndiff >>
rect 70 489 100 500
rect 70 471 76 489
rect 94 471 100 489
rect 70 453 100 471
rect 70 435 76 453
rect 94 435 100 453
rect 70 417 100 435
rect 70 399 76 417
rect 94 399 100 417
rect 70 381 100 399
rect 70 363 76 381
rect 94 363 100 381
rect 70 345 100 363
rect 70 327 76 345
rect 94 327 100 345
rect 70 309 100 327
rect 70 291 76 309
rect 94 291 100 309
rect 70 273 100 291
rect 70 255 76 273
rect 94 255 100 273
rect 70 237 100 255
rect 70 219 76 237
rect 94 219 100 237
rect 70 201 100 219
rect 70 183 76 201
rect 94 183 100 201
rect 70 165 100 183
rect 70 147 76 165
rect 94 147 100 165
rect 70 129 100 147
rect 70 111 76 129
rect 94 111 100 129
rect 70 93 100 111
rect 70 75 76 93
rect 94 75 100 93
rect 70 57 100 75
rect 70 39 76 57
rect 94 39 100 57
rect 70 21 100 39
rect 70 3 76 21
rect 94 3 100 21
rect 70 -15 100 3
rect 70 -33 76 -15
rect 94 -33 100 -15
rect 70 -51 100 -33
rect 70 -69 76 -51
rect 94 -69 100 -51
rect 70 -100 100 -69
rect 450 489 480 500
rect 450 471 456 489
rect 474 471 480 489
rect 450 453 480 471
rect 450 435 456 453
rect 474 435 480 453
rect 450 417 480 435
rect 450 399 456 417
rect 474 399 480 417
rect 450 381 480 399
rect 450 363 456 381
rect 474 363 480 381
rect 450 345 480 363
rect 450 327 456 345
rect 474 327 480 345
rect 450 309 480 327
rect 450 291 456 309
rect 474 291 480 309
rect 450 273 480 291
rect 450 255 456 273
rect 474 255 480 273
rect 450 237 480 255
rect 450 219 456 237
rect 474 219 480 237
rect 450 201 480 219
rect 450 183 456 201
rect 474 183 480 201
rect 450 165 480 183
rect 450 147 456 165
rect 474 147 480 165
rect 450 129 480 147
rect 450 111 456 129
rect 474 111 480 129
rect 450 93 480 111
rect 450 75 456 93
rect 474 75 480 93
rect 450 57 480 75
rect 450 39 456 57
rect 474 39 480 57
rect 450 21 480 39
rect 450 3 456 21
rect 474 3 480 21
rect 450 -15 480 3
rect 450 -33 456 -15
rect 474 -33 480 -15
rect 450 -51 480 -33
rect 450 -69 456 -51
rect 474 -69 480 -51
rect 450 -100 480 -69
<< ndiffc >>
rect 76 471 94 489
rect 76 435 94 453
rect 76 399 94 417
rect 76 363 94 381
rect 76 327 94 345
rect 76 291 94 309
rect 76 255 94 273
rect 76 219 94 237
rect 76 183 94 201
rect 76 147 94 165
rect 76 111 94 129
rect 76 75 94 93
rect 76 39 94 57
rect 76 3 94 21
rect 76 -33 94 -15
rect 76 -69 94 -51
rect 456 471 474 489
rect 456 435 474 453
rect 456 399 474 417
rect 456 363 474 381
rect 456 327 474 345
rect 456 291 474 309
rect 456 255 474 273
rect 456 219 474 237
rect 456 183 474 201
rect 456 147 474 165
rect 456 111 474 129
rect 456 75 474 93
rect 456 39 474 57
rect 456 3 474 21
rect 456 -33 474 -15
rect 456 -69 474 -51
<< poly >>
rect 100 500 450 520
rect 100 -120 450 -100
<< locali >>
rect 70 489 100 502
rect 70 471 76 489
rect 94 471 100 489
rect 70 453 100 471
rect 70 435 76 453
rect 94 435 100 453
rect 70 417 100 435
rect 70 399 76 417
rect 94 399 100 417
rect 70 381 100 399
rect 70 363 76 381
rect 94 363 100 381
rect 70 345 100 363
rect 70 327 76 345
rect 94 327 100 345
rect 70 309 100 327
rect 70 291 76 309
rect 94 291 100 309
rect 70 273 100 291
rect 70 255 76 273
rect 94 255 100 273
rect 70 237 100 255
rect 70 219 76 237
rect 94 219 100 237
rect 70 201 100 219
rect 70 183 76 201
rect 94 183 100 201
rect 70 165 100 183
rect 70 147 76 165
rect 94 147 100 165
rect 70 129 100 147
rect 70 111 76 129
rect 94 111 100 129
rect 70 93 100 111
rect 70 75 76 93
rect 94 75 100 93
rect 70 57 100 75
rect 70 39 76 57
rect 94 39 100 57
rect 70 21 100 39
rect 70 3 76 21
rect 94 3 100 21
rect 70 -15 100 3
rect 70 -33 76 -15
rect 94 -33 100 -15
rect 70 -51 100 -33
rect 70 -69 76 -51
rect 94 -69 100 -51
rect 70 -102 100 -69
rect 450 489 480 502
rect 450 471 456 489
rect 474 471 480 489
rect 450 453 480 471
rect 450 435 456 453
rect 474 435 480 453
rect 450 417 480 435
rect 450 399 456 417
rect 474 399 480 417
rect 450 381 480 399
rect 450 363 456 381
rect 474 363 480 381
rect 450 345 480 363
rect 450 327 456 345
rect 474 327 480 345
rect 450 309 480 327
rect 450 291 456 309
rect 474 291 480 309
rect 450 273 480 291
rect 450 255 456 273
rect 474 255 480 273
rect 450 237 480 255
rect 450 219 456 237
rect 474 219 480 237
rect 450 201 480 219
rect 450 183 456 201
rect 474 183 480 201
rect 450 165 480 183
rect 450 147 456 165
rect 474 147 480 165
rect 450 129 480 147
rect 450 111 456 129
rect 474 111 480 129
rect 450 93 480 111
rect 450 75 456 93
rect 474 75 480 93
rect 450 57 480 75
rect 450 39 456 57
rect 474 39 480 57
rect 450 21 480 39
rect 450 3 456 21
rect 474 3 480 21
rect 450 -15 480 3
rect 450 -33 456 -15
rect 474 -33 480 -15
rect 450 -51 480 -33
rect 450 -69 456 -51
rect 474 -69 480 -51
rect 450 -102 480 -69
<< labels >>
rlabel locali 85 500 85 500 1 D
rlabel locali 465 500 465 500 1 S
rlabel pwell 480 520 480 520 1 B
rlabel poly 270 510 270 510 1 G
<< end >>
