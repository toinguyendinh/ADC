* NGSPICE file created from main_inv.ext - technology: sky130A

.subckt main_inv A VPWR VGND Y
X0 VPWR A Y VDD sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.3 ps=2.3 w=2 l=0.5
X1 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.3 ps=2.6 w=1 l=0.5
X2 VGND A Y GND sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.15 ps=1.3 w=1 l=0.5
X3 Y A VGND GND sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.5
X4 Y A VPWR VDD sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.3 ps=2.3 w=2 l=0.5
X5 Y A VPWR VDD sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.6 ps=4.6 w=2 l=0.5
X6 VPWR A Y VDD sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.3 ps=2.3 w=2 l=0.5
X7 VGND A Y GND sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.15 ps=1.3 w=1 l=0.5
.ends

