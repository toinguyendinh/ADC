magic
tech sky130A
timestamp 1692022408
<< pwell >>
rect -50 -40 400 360
<< nmos >>
rect 0 0 350 320
<< ndiff >>
rect -30 309 0 320
rect -30 291 -24 309
rect -6 291 0 309
rect -30 273 0 291
rect -30 255 -24 273
rect -6 255 0 273
rect -30 237 0 255
rect -30 219 -24 237
rect -6 219 0 237
rect -30 201 0 219
rect -30 183 -24 201
rect -6 183 0 201
rect -30 165 0 183
rect -30 147 -24 165
rect -6 147 0 165
rect -30 129 0 147
rect -30 111 -24 129
rect -6 111 0 129
rect -30 93 0 111
rect -30 75 -24 93
rect -6 75 0 93
rect -30 57 0 75
rect -30 39 -24 57
rect -6 39 0 57
rect -30 0 0 39
rect 350 309 380 320
rect 350 291 356 309
rect 374 291 380 309
rect 350 273 380 291
rect 350 255 356 273
rect 374 255 380 273
rect 350 237 380 255
rect 350 219 356 237
rect 374 219 380 237
rect 350 201 380 219
rect 350 183 356 201
rect 374 183 380 201
rect 350 165 380 183
rect 350 147 356 165
rect 374 147 380 165
rect 350 129 380 147
rect 350 111 356 129
rect 374 111 380 129
rect 350 93 380 111
rect 350 75 356 93
rect 374 75 380 93
rect 350 57 380 75
rect 350 39 356 57
rect 374 39 380 57
rect 350 0 380 39
<< ndiffc >>
rect -24 291 -6 309
rect -24 255 -6 273
rect -24 219 -6 237
rect -24 183 -6 201
rect -24 147 -6 165
rect -24 111 -6 129
rect -24 75 -6 93
rect -24 39 -6 57
rect 356 291 374 309
rect 356 255 374 273
rect 356 219 374 237
rect 356 183 374 201
rect 356 147 374 165
rect 356 111 374 129
rect 356 75 374 93
rect 356 39 374 57
<< poly >>
rect 0 320 350 340
rect 0 -20 350 0
<< locali >>
rect -30 309 0 322
rect -30 291 -24 309
rect -6 291 0 309
rect -30 273 0 291
rect -30 255 -24 273
rect -6 255 0 273
rect -30 237 0 255
rect -30 219 -24 237
rect -6 219 0 237
rect -30 201 0 219
rect -30 183 -24 201
rect -6 183 0 201
rect -30 165 0 183
rect -30 147 -24 165
rect -6 147 0 165
rect -30 129 0 147
rect -30 111 -24 129
rect -6 111 0 129
rect -30 93 0 111
rect -30 75 -24 93
rect -6 75 0 93
rect -30 57 0 75
rect -30 39 -24 57
rect -6 39 0 57
rect -30 -2 0 39
rect 350 309 380 322
rect 350 291 356 309
rect 374 291 380 309
rect 350 273 380 291
rect 350 255 356 273
rect 374 255 380 273
rect 350 237 380 255
rect 350 219 356 237
rect 374 219 380 237
rect 350 201 380 219
rect 350 183 356 201
rect 374 183 380 201
rect 350 165 380 183
rect 350 147 356 165
rect 374 147 380 165
rect 350 129 380 147
rect 350 111 356 129
rect 374 111 380 129
rect 350 93 380 111
rect 350 75 356 93
rect 374 75 380 93
rect 350 57 380 75
rect 350 39 356 57
rect 374 39 380 57
rect 350 -2 380 39
<< labels >>
rlabel locali -15 320 -15 320 1 D
rlabel locali 365 322 365 322 1 S
rlabel poly 170 330 170 330 1 G
rlabel pwell 380 340 380 340 1 B
<< end >>
