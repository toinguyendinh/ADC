magic
tech sky130A
timestamp 1699711427
<< nwell >>
rect -50 150 390 410
<< pwell >>
rect -50 -4 390 130
rect -50 -20 50 -4
rect 80 -20 210 -4
rect 240 -20 390 -4
rect -50 -30 390 -20
rect 350 -50 370 -30
<< nmos >>
rect 0 0 50 100
rect 80 0 130 100
rect 160 0 210 100
rect 240 0 290 100
<< pmos >>
rect 0 180 50 380
rect 80 180 130 380
rect 160 180 210 380
rect 240 180 290 380
<< ndiff >>
rect -30 96 0 100
rect -30 78 -24 96
rect -6 78 0 96
rect -30 60 0 78
rect -30 40 -24 60
rect -6 40 0 60
rect -30 22 0 40
rect -30 4 -24 22
rect -6 4 0 22
rect -30 0 0 4
rect 50 96 80 100
rect 50 78 56 96
rect 74 78 80 96
rect 50 60 80 78
rect 50 40 56 60
rect 74 40 80 60
rect 50 22 80 40
rect 50 4 56 22
rect 74 4 80 22
rect 50 0 80 4
rect 130 96 160 100
rect 130 78 136 96
rect 154 78 160 96
rect 130 60 160 78
rect 130 40 136 60
rect 154 40 160 60
rect 130 22 160 40
rect 130 4 136 22
rect 154 4 160 22
rect 130 0 160 4
rect 210 96 240 100
rect 210 78 216 96
rect 234 78 240 96
rect 210 60 240 78
rect 210 40 216 60
rect 234 40 240 60
rect 210 22 240 40
rect 210 4 216 22
rect 234 4 240 22
rect 210 0 240 4
rect 290 96 320 100
rect 290 78 296 96
rect 314 78 320 96
rect 290 60 320 78
rect 290 40 296 60
rect 314 40 320 60
rect 290 22 320 40
rect 290 4 296 22
rect 314 4 320 22
rect 290 0 320 4
<< pdiff >>
rect -30 376 0 380
rect -30 358 -24 376
rect -6 358 0 376
rect -30 340 0 358
rect -30 320 -24 340
rect -6 320 0 340
rect -30 302 0 320
rect -30 258 -24 302
rect -6 258 0 302
rect -30 240 0 258
rect -30 220 -24 240
rect -6 220 0 240
rect -30 202 0 220
rect -30 184 -24 202
rect -6 184 0 202
rect -30 180 0 184
rect 50 376 80 380
rect 50 358 56 376
rect 74 358 80 376
rect 50 340 80 358
rect 50 320 56 340
rect 74 320 80 340
rect 50 302 80 320
rect 50 258 56 302
rect 74 258 80 302
rect 50 240 80 258
rect 50 220 56 240
rect 74 220 80 240
rect 50 202 80 220
rect 50 184 56 202
rect 74 184 80 202
rect 50 180 80 184
rect 130 376 160 380
rect 130 358 136 376
rect 154 358 160 376
rect 130 340 160 358
rect 130 320 136 340
rect 154 320 160 340
rect 130 302 160 320
rect 130 258 136 302
rect 154 258 160 302
rect 130 240 160 258
rect 130 220 136 240
rect 154 220 160 240
rect 130 202 160 220
rect 130 184 136 202
rect 154 184 160 202
rect 130 180 160 184
rect 210 376 240 380
rect 210 358 216 376
rect 234 358 240 376
rect 210 340 240 358
rect 210 320 216 340
rect 234 320 240 340
rect 210 302 240 320
rect 210 258 216 302
rect 234 258 240 302
rect 210 240 240 258
rect 210 220 216 240
rect 234 220 240 240
rect 210 202 240 220
rect 210 184 216 202
rect 234 184 240 202
rect 210 180 240 184
rect 290 376 320 380
rect 290 358 296 376
rect 314 358 320 376
rect 290 340 320 358
rect 290 320 296 340
rect 314 320 320 340
rect 290 302 320 320
rect 290 258 296 302
rect 314 258 320 302
rect 290 240 320 258
rect 290 220 296 240
rect 314 220 320 240
rect 290 202 320 220
rect 290 184 296 202
rect 314 184 320 202
rect 290 180 320 184
<< ndiffc >>
rect -24 78 -6 96
rect -24 40 -6 60
rect -24 4 -6 22
rect 56 78 74 96
rect 56 40 74 60
rect 56 4 74 22
rect 136 78 154 96
rect 136 40 154 60
rect 136 4 154 22
rect 216 78 234 96
rect 216 40 234 60
rect 216 4 234 22
rect 296 78 314 96
rect 296 40 314 60
rect 296 4 314 22
<< pdiffc >>
rect -24 358 -6 376
rect -24 320 -6 340
rect -24 258 -6 302
rect -24 220 -6 240
rect -24 184 -6 202
rect 56 358 74 376
rect 56 320 74 340
rect 56 258 74 302
rect 56 220 74 240
rect 56 184 74 202
rect 136 358 154 376
rect 136 320 154 340
rect 136 258 154 302
rect 136 220 154 240
rect 136 184 154 202
rect 216 358 234 376
rect 216 320 234 340
rect 216 258 234 302
rect 216 220 234 240
rect 216 184 234 202
rect 296 358 314 376
rect 296 320 314 340
rect 296 258 314 302
rect 296 220 314 240
rect 296 184 314 202
<< psubdiff >>
rect 350 96 370 112
rect 350 60 370 78
rect 350 22 370 40
rect 350 -12 370 4
<< nsubdiff >>
rect 350 376 370 392
rect 350 340 370 358
rect 350 302 370 320
rect 350 240 370 258
rect 350 202 370 220
rect 350 168 370 184
<< psubdiffcont >>
rect 350 78 370 96
rect 350 40 370 60
rect 350 4 370 22
<< nsubdiffcont >>
rect 350 358 370 376
rect 350 320 370 340
rect 350 258 370 302
rect 350 220 370 240
rect 350 184 370 202
<< poly >>
rect 0 380 50 400
rect 80 380 130 400
rect 160 380 210 400
rect 240 380 290 400
rect 0 160 50 180
rect 80 160 130 180
rect 160 160 210 180
rect 240 160 290 180
rect 0 120 290 160
rect 0 100 50 120
rect 80 100 130 120
rect 160 100 210 120
rect 240 100 290 120
rect 0 -20 50 0
rect 80 -20 130 0
rect 160 -20 210 0
rect 240 -20 290 0
<< locali >>
rect -30 410 320 430
rect -30 376 0 410
rect -30 358 -24 376
rect -6 358 0 376
rect -30 340 0 358
rect -30 320 -24 340
rect -6 320 0 340
rect -30 302 0 320
rect -30 258 -24 302
rect -6 258 0 302
rect -30 240 0 258
rect -30 220 -24 240
rect -6 220 0 240
rect -30 202 0 220
rect -30 184 -24 202
rect -6 184 0 202
rect -30 176 0 184
rect 50 376 80 384
rect 50 358 56 376
rect 74 358 80 376
rect 50 340 80 358
rect 50 320 56 340
rect 74 320 80 340
rect 50 302 80 320
rect 50 258 56 302
rect 74 258 80 302
rect 50 240 80 258
rect 50 220 56 240
rect 74 220 80 240
rect 50 202 80 220
rect 50 184 56 202
rect 74 184 80 202
rect 50 155 80 184
rect 130 376 160 410
rect 130 358 136 376
rect 154 358 160 376
rect 130 340 160 358
rect 130 320 136 340
rect 154 320 160 340
rect 130 302 160 320
rect 130 258 136 302
rect 154 258 160 302
rect 130 240 160 258
rect 130 220 136 240
rect 154 220 160 240
rect 130 202 160 220
rect 130 184 136 202
rect 154 184 160 202
rect 130 176 160 184
rect 210 376 240 384
rect 210 358 216 376
rect 234 358 240 376
rect 210 340 240 358
rect 210 320 216 340
rect 234 320 240 340
rect 210 302 240 320
rect 210 258 216 302
rect 234 258 240 302
rect 210 240 240 258
rect 210 220 216 240
rect 234 220 240 240
rect 210 202 240 220
rect 210 184 216 202
rect 234 184 240 202
rect 210 155 240 184
rect 290 376 320 410
rect 290 358 296 376
rect 314 358 320 376
rect 290 340 320 358
rect 290 320 296 340
rect 314 320 320 340
rect 290 302 320 320
rect 290 258 296 302
rect 314 258 320 302
rect 290 240 320 258
rect 290 220 296 240
rect 314 220 320 240
rect 290 202 320 220
rect 290 184 296 202
rect 314 184 320 202
rect 290 176 320 184
rect 350 376 370 430
rect 350 340 370 358
rect 350 302 370 320
rect 350 240 370 258
rect 350 202 370 220
rect 350 172 370 184
rect 50 125 370 155
rect -30 96 0 104
rect -30 78 -24 96
rect -6 78 0 96
rect -30 60 0 78
rect -30 40 -24 60
rect -6 40 0 60
rect -30 22 0 40
rect -30 4 -24 22
rect -6 4 0 22
rect -30 -30 0 4
rect 50 96 80 125
rect 50 78 56 96
rect 74 78 80 96
rect 50 60 80 78
rect 50 40 56 60
rect 74 40 80 60
rect 50 22 80 40
rect 50 4 56 22
rect 74 4 80 22
rect 50 -4 80 4
rect 130 96 160 104
rect 130 78 136 96
rect 154 78 160 96
rect 130 60 160 78
rect 130 40 136 60
rect 154 40 160 60
rect 130 22 160 40
rect 130 4 136 22
rect 154 4 160 22
rect 130 -30 160 4
rect 210 96 240 125
rect 210 78 216 96
rect 234 78 240 96
rect 210 60 240 78
rect 210 40 216 60
rect 234 40 240 60
rect 210 22 240 40
rect 210 4 216 22
rect 234 4 240 22
rect 210 -4 240 4
rect 290 96 320 104
rect 290 78 296 96
rect 314 78 320 96
rect 290 60 320 78
rect 290 40 296 60
rect 314 40 320 60
rect 290 22 320 40
rect 290 4 296 22
rect 314 4 320 22
rect 290 -30 320 4
rect -30 -50 320 -30
rect 350 96 370 108
rect 350 60 370 78
rect 350 22 370 40
rect 350 -50 370 4
<< labels >>
rlabel poly 0 140 0 140 1 A
port 1 n default input
rlabel locali -30 400 -30 400 1 VPWR
port 2 n
rlabel locali -30 -20 -30 -20 1 VGND
port 3 n
rlabel locali 360 -45 360 -45 1 GND
rlabel locali 370 140 370 140 1 Y
port 4 n
rlabel locali 360 425 360 425 5 VDD
<< end >>
