**.subckt NMOS
VG G GND 0
VD D GND 0
XM1 D G GND 0 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
**** begin user architecture code


.lib /home/dkits/efabless/mpw-5/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.inc /home/dkits/efabless/mpw-5/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice




.control
set nobreak
set numthread=11

dc VD 0 2 0.01 VG 0 2 0.2
print format=raw file=NMOS.raw v(*) i(*)

.endc


**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes
.end
