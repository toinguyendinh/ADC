magic
tech sky130A
timestamp 1692027968
<< nwell >>
rect 0 0 450 680
<< pmos >>
rect 50 40 400 640
<< pdiff >>
rect 20 629 50 640
rect 20 611 26 629
rect 44 611 50 629
rect 20 593 50 611
rect 20 575 26 593
rect 44 575 50 593
rect 20 557 50 575
rect 20 539 26 557
rect 44 539 50 557
rect 20 521 50 539
rect 20 503 26 521
rect 44 503 50 521
rect 20 485 50 503
rect 20 467 26 485
rect 44 467 50 485
rect 20 449 50 467
rect 20 431 26 449
rect 44 431 50 449
rect 20 413 50 431
rect 20 395 26 413
rect 44 395 50 413
rect 20 377 50 395
rect 20 359 26 377
rect 44 359 50 377
rect 20 341 50 359
rect 20 323 26 341
rect 44 323 50 341
rect 20 305 50 323
rect 20 287 26 305
rect 44 287 50 305
rect 20 269 50 287
rect 20 251 26 269
rect 44 251 50 269
rect 20 233 50 251
rect 20 215 26 233
rect 44 215 50 233
rect 20 197 50 215
rect 20 179 26 197
rect 44 179 50 197
rect 20 161 50 179
rect 20 143 26 161
rect 44 143 50 161
rect 20 125 50 143
rect 20 107 26 125
rect 44 107 50 125
rect 20 89 50 107
rect 20 71 26 89
rect 44 71 50 89
rect 20 40 50 71
rect 400 629 430 640
rect 400 611 406 629
rect 424 611 430 629
rect 400 593 430 611
rect 400 575 406 593
rect 424 575 430 593
rect 400 557 430 575
rect 400 539 406 557
rect 424 539 430 557
rect 400 521 430 539
rect 400 503 406 521
rect 424 503 430 521
rect 400 485 430 503
rect 400 467 406 485
rect 424 467 430 485
rect 400 449 430 467
rect 400 431 406 449
rect 424 431 430 449
rect 400 413 430 431
rect 400 395 406 413
rect 424 395 430 413
rect 400 377 430 395
rect 400 359 406 377
rect 424 359 430 377
rect 400 341 430 359
rect 400 323 406 341
rect 424 323 430 341
rect 400 305 430 323
rect 400 287 406 305
rect 424 287 430 305
rect 400 269 430 287
rect 400 251 406 269
rect 424 251 430 269
rect 400 233 430 251
rect 400 215 406 233
rect 424 215 430 233
rect 400 197 430 215
rect 400 179 406 197
rect 424 179 430 197
rect 400 161 430 179
rect 400 143 406 161
rect 424 143 430 161
rect 400 125 430 143
rect 400 107 406 125
rect 424 107 430 125
rect 400 89 430 107
rect 400 71 406 89
rect 424 71 430 89
rect 400 40 430 71
<< pdiffc >>
rect 26 611 44 629
rect 26 575 44 593
rect 26 539 44 557
rect 26 503 44 521
rect 26 467 44 485
rect 26 431 44 449
rect 26 395 44 413
rect 26 359 44 377
rect 26 323 44 341
rect 26 287 44 305
rect 26 251 44 269
rect 26 215 44 233
rect 26 179 44 197
rect 26 143 44 161
rect 26 107 44 125
rect 26 71 44 89
rect 406 611 424 629
rect 406 575 424 593
rect 406 539 424 557
rect 406 503 424 521
rect 406 467 424 485
rect 406 431 424 449
rect 406 395 424 413
rect 406 359 424 377
rect 406 323 424 341
rect 406 287 424 305
rect 406 251 424 269
rect 406 215 424 233
rect 406 179 424 197
rect 406 143 424 161
rect 406 107 424 125
rect 406 71 424 89
<< poly >>
rect 50 640 400 660
rect 50 20 400 40
<< locali >>
rect 20 629 50 642
rect 20 611 26 629
rect 44 611 50 629
rect 20 593 50 611
rect 20 575 26 593
rect 44 575 50 593
rect 20 557 50 575
rect 20 539 26 557
rect 44 539 50 557
rect 20 521 50 539
rect 20 503 26 521
rect 44 503 50 521
rect 20 485 50 503
rect 20 467 26 485
rect 44 467 50 485
rect 20 449 50 467
rect 20 431 26 449
rect 44 431 50 449
rect 20 413 50 431
rect 20 395 26 413
rect 44 395 50 413
rect 20 377 50 395
rect 20 359 26 377
rect 44 359 50 377
rect 20 341 50 359
rect 20 323 26 341
rect 44 323 50 341
rect 20 305 50 323
rect 20 287 26 305
rect 44 287 50 305
rect 20 269 50 287
rect 20 251 26 269
rect 44 251 50 269
rect 20 233 50 251
rect 20 215 26 233
rect 44 215 50 233
rect 20 197 50 215
rect 20 179 26 197
rect 44 179 50 197
rect 20 161 50 179
rect 20 143 26 161
rect 44 143 50 161
rect 20 125 50 143
rect 20 107 26 125
rect 44 107 50 125
rect 20 89 50 107
rect 20 71 26 89
rect 44 71 50 89
rect 20 38 50 71
rect 400 629 430 642
rect 400 611 406 629
rect 424 611 430 629
rect 400 593 430 611
rect 400 575 406 593
rect 424 575 430 593
rect 400 557 430 575
rect 400 539 406 557
rect 424 539 430 557
rect 400 521 430 539
rect 400 503 406 521
rect 424 503 430 521
rect 400 485 430 503
rect 400 467 406 485
rect 424 467 430 485
rect 400 449 430 467
rect 400 431 406 449
rect 424 431 430 449
rect 400 413 430 431
rect 400 395 406 413
rect 424 395 430 413
rect 400 377 430 395
rect 400 359 406 377
rect 424 359 430 377
rect 400 341 430 359
rect 400 323 406 341
rect 424 323 430 341
rect 400 305 430 323
rect 400 287 406 305
rect 424 287 430 305
rect 400 269 430 287
rect 400 251 406 269
rect 424 251 430 269
rect 400 233 430 251
rect 400 215 406 233
rect 424 215 430 233
rect 400 197 430 215
rect 400 179 406 197
rect 424 179 430 197
rect 400 161 430 179
rect 400 143 406 161
rect 424 143 430 161
rect 400 125 430 143
rect 400 107 406 125
rect 424 107 430 125
rect 400 89 430 107
rect 400 71 406 89
rect 424 71 430 89
rect 400 38 430 71
<< labels >>
rlabel locali 35 40 35 40 1 D
rlabel poly 220 40 220 40 1 G
rlabel locali 415 40 415 40 1 S
rlabel nwell 430 20 430 20 1 B
<< end >>
